magic
tech sky130A
timestamp 1756722359
<< locali >>
rect -48 -1251 48 -1118
rect 527 -1251 623 -1120
rect -48 -1253 623 -1251
rect -48 -1343 147 -1253
rect 237 -1343 623 -1253
rect -48 -1347 623 -1343
<< viali >>
rect 147 -1343 237 -1253
<< metal1 >>
rect 80 -41 112 458
rect 77 -73 80 -41
rect 112 -73 115 -41
rect 80 -857 112 -73
rect 144 -1253 240 745
rect 336 644 600 740
rect 504 333 600 644
rect 336 237 600 333
rect 389 -41 421 -38
rect 389 -76 421 -73
rect 504 -452 600 237
rect 336 -548 600 -452
rect 504 -954 600 -548
rect 337 -1050 600 -954
rect 144 -1343 147 -1253
rect 237 -1343 240 -1253
rect 144 -1349 240 -1343
<< via1 >>
rect 80 -73 112 -41
rect 389 -73 421 -41
<< metal2 >>
rect 80 -41 112 -38
rect -90 -73 80 -41
rect 112 -73 389 -41
rect 421 -73 424 -41
rect 80 -76 112 -73
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1756722359
transform 1 0 0 0 1 401
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1756722359
transform 1 0 0 0 1 -1203
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1756722359
transform 1 0 0 0 1 0
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1756722359
transform 1 0 0 0 1 -400
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1756722359
transform 1 0 0 0 1 -799
box -92 -64 668 464
<< labels >>
flabel locali -42 -1347 54 -1251 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel metal1 513 -1027 576 696 0 FreeSans 800 0 0 0 IBNS_20U
port 0 nsew
flabel metal2 -88 -72 69 -44 0 FreeSans 800 0 0 0 IBPS_5U
port 2 nsew
<< end >>
